// PLACEHOLDER FOR ENV SETUP

module rt_ss_wrapper_0 #()();


rt_top #() i_rt_top ();

endmodule : rt_ss_wrapper_0